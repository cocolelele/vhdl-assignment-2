
entity jkhgvkjhg is
    Port ( X : in  BIT_VECTOR (7 downto 0);
           Y : in  BIT_VECTOR (7 downto 0);
           Start : in  BIT;
           CLK : in  BIT;
           Reset : in  BIT;
           Result : out  BIT_VECTOR (15 downto 0);
           Done : out  BIT);
end jkhgvkjhg;

architecture Behavioral of jkhgvkjhg is

begin


end Behavioral;

